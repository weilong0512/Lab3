savavs